`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:49:07 05/09/2017 
// Design Name: 
// Module Name:    Shifter_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Shifter_2(
    input [31:0] Input,
    output [31:0] Output
    );
	 
	 assign Output = Input ;


endmodule
