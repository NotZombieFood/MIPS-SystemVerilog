��` t i m e s c a l e   1 n s   /   1 p s  
 / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / /  
 / /   C o m p a n y :    
 / /   E n g i n e e r :    
 / /    
 / /   C r e a t e   D a t e :         2 2 : 0 3 : 2 0   0 5 / 0 9 / 2 0 1 7    
 / /   D e s i g n   N a m e :    
 / /   M o d u l e   N a m e :         P C    
 / /   P r o j e c t   N a m e :    
 / /   T a r g e t   D e v i c e s :    
 / /   T o o l   v e r s i o n s :    
 / /   D e s c r i p t i o n :    
 / /  
 / /   D e p e n d e n c i e s :    
 / /  
 / /   R e v i s i o n :    
 / /   R e v i s i o n   0 . 0 1   -   F i l e   C r e a t e d  
 / /   A d d i t i o n a l   C o m m e n t s :    
 / /  
 / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / /  
 m o d u l e   I n s t r u c t i o n M e m o r y (  
         i n p u t   [ 3 1 : 0 ]   A d d r e s s ,  
         o u t p u t   l o g i c   [ 3 1 : 0 ]   W o r d  
         ) ;  
 / / u s e   6   b i t s   f o r   a d r e s s 	  
 a l w a y s _ c o m b   b e g i n  
 	 c a s e   ( A d d r e s s [ 7 : 0 ] )  
 	 	 	 0 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 - 0 1 0 0 1 0 0 0 ;   	 / / I n s t r u c t i o n   0 *  
 	 	 	 4 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 - 0 1 0 0 0 1 0 1 ; 	 	 / / I n s t r u c t i o n   4 *  
 	 	 	 8 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 - - 0 1 0 0 1 1 0 0 ; 	 	 / / I n s t r u c t i o n   8 *  
 	 	 	 1 2 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 - - 0 1 0 0 1 1 0 0 ;   	 / / I n s t r u c t i o n   1 2 *  
 	 	 	 1 6 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 - 0 1 0 0 1 1 1 1 ;   	 / / I n s t r u c t i o n   1 6 *  
 	 	 	 2 0 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 - - 0 0 1 0 0 0 0 0 , , , ;   	 / / I n s t r u c t i o n   2 0 *  
 	 	 	 2 4 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 - 0 1 0 1 0 1 1 1 ;   	 / / I n s t r u c t i o n   2 4 *  
 	 	 	 2 8 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 - 0 1 0 0 1 1 1 1 ;   	 / / I n s t r u c t i o n   2 8 *  
 	 	 	 3 2 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 - - 0 1 0 1 0 0 1 0 , ;   	 / / I n s t r u c t i o n   3 2 *  
 	 	 	 3 6 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 - - 0 1 0 0 1 1 0 0 ;   	 / / I n s t r u c t i o n   3 6 *  
 	 	 	 4 0 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 - - - 0 1 0 0 0 1 0 0 ;   	 / / I n s t r u c t i o n   4 0 *  
 	 	 	 4 4 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 , 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ;   	 / / I n s t r u c t i o n   4 4 *  
 	 	 	 4 8 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 ;   	 / / I n s t r u c t i o n   4 8 *  
 	 	 	 5 2 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 ;   	 / / I n s t r u c t i o n   5 2 *  
 	 	 	 5 6 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 ;   	 / / I n s t r u c t i o n   5 6 *  
 	 	 	 6 0 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 ;   	 / / I n s t r u c t i o n   6 0 *  
 	 	 	 6 4 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 ;   	 / / I n s t r u c t i o n   6 4 *  
 	 	 	 6 8 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 ;   	 / / I n s t r u c t i o n   6 8 *  
 	 	 	 7 2 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 ;   	 / / I n s t r u c t i o n   7 2 *  
 	 	 	 7 6 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 ;   	 / / I n s t r u c t i o n   7 6 *  
 	 	 	 8 0 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 , 0 0 0 0 0 , 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 ;   	 / / I n s t r u c t i o n   8 0 *  
 	 	 	 8 4 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 ;   	 / / I n s t r u c t i o n   8 4 *  
 	 	 	 8 8 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 ;   	 / / I n s t r u c t i o n   8 8 *  
 	 	 	 9 2 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 ;   	 / / I n s t r u c t i o n   9 2 *  
 	 	 	 9 6 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 , 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 ;   	 / / I n s t r u c t i o n   9 6 *  
 	 	 	 1 0 0 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 , 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 ;   	 / / I n s t r u c t i o n   1 0 0 *  
 	 	 	 1 0 4 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 - 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 ;   	 / / I n s t r u c t i o n   1 0 4 *  
 	 	 	 1 0 8 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 ;   	 / / I n s t r u c t i o n   1 0 8 *  
 	 	 	 1 1 2 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 , 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 ;   	 / / I n s t r u c t i o n   1 1 2 *  
 	 	 	 1 1 6 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 ;   	 / / I n s t r u c t i o n   1 1 6 *  
 	 	 	 1 2 0 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 , 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 ;   	 / / I n s t r u c t i o n   1 2 0 *  
 	 	 	 1 2 4 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 ;   	 / / I n s t r u c t i o n   1 2 4 *  
 	 	 	 1 2 8 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 ;   	 / / I n s t r u c t i o n   1 2 8 *  
 	 	 	 1 3 2 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 ;   	 / / I n s t r u c t i o n   1 3 2  
 	 	 	 1 3 6 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 ; 	 / / I n s t r u c t i o n   1 3 6 *  
 	 	 	 1 4 0 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 ; 	 / / I n s t r u c t i o n   1 4 0 *  
 	 	 	 1 4 4 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 , 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 ; 	 / / I n s t r u c t i o n   1 4 4 *  
 	 	 	 1 4 8 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 ; 	 / / I n s t r u c t i o n   1 4 8 *  
 	 	 	 1 5 2 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 ; 	 / / I n s t r u c t i o n   1 5 2 *  
 	 	 	 1 5 6 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 1 ; 	 / / I n s t r u c t i o n   1 5 6 *  
 	 	 	 1 6 0 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 , 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 ; 	 / / I n s t r u c t i o n   1 6 0 *  
 	 	 	 1 6 4 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 ; 	 / / I n s t r u c t i o n   1 6 4 *  
 	 	 	 1 6 8 :   W o r d   =   3 2 ' b 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ; 	 / / I n s t r u c t i o n   1 6 8 *  
 	 	 	 1 7 2 :   W o r d   =   3 2 ' b 1 0 1 0 1 1 0 0 0 0 0 , 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 ; 	 / / I n s t r u c t i o n   1 7 2 *  
 	 	 	 1 7 6 :   W o r d   =   3 2 ' b 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 - 1 0 1 1 0 0 0 0 , ; 	 / / I n s t r u c t i o n   1 7 6 *  
 	 	 	 d e f a u l t :   W o r d   =   3 2 ' b 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ;  
 	 e n d c a s e    
 e n d  
 e n d m o d u l e  
 